CIRCUIT C:\microwind2\Book on CMOS\AmpliDiffNP.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
VVp 9 0 PULSE(0.00 1.20 2.00N 14.00N 14.00N 2.00N 32.00N)
V10_Vbias 10 0 DC 0.60V
V11_VbiasP 11 0 DC 0.60V
*
* List of nodes
* "Vout" corresponds to n�3
* "N4" corresponds to n�4
* "nMOS current mirror" corresponds to n�5
* "pMOS current mirror" corresponds to n�7
* "N8" corresponds to n�8
* "Vp" corresponds to n�9
* "Vbias" corresponds to n�10
* "VbiasP" corresponds to n�11
*
* MOS devices
MN1 0 5 3 0 N1  W= 0.84U L= 0.60U
MN2 5 5 0 0 N1  W= 0.84U L= 0.60U
MN3 8 3 3 0 N1  W= 0.54U L= 0.60U
MN4 7 9 8 0 N1  W= 0.54U L= 0.60U
MN5 0 10 8 0 N1  W= 0.54U L= 0.60U
MP1 4 3 3 1 P1  W= 0.54U L= 0.60U
MP2 5 9 4 1 P1  W= 0.54U L= 0.60U
MP3 1 11 4 1 P1  W= 0.54U L= 0.60U
MP4 1 7 3 1 P1  W= 0.84U L= 0.60U
MP5 7 7 1 1 P1  W= 0.84U L= 0.60U
*
C2 1 0  7.333fF
C3 3 0  1.855fF
C4 4 0  0.442fF
C5 5 0  1.330fF
C7 7 0  1.325fF
C8 8 0  0.501fF
C9 9 0  0.890fF
C10 10 0  0.337fF
C11 11 0  0.337fF
*
*
* n-MOS BSIM4 :
* low leakage
.MODEL N1 NMOS LEVEL=14 VTO=0.40 U0=0.050 TOX= 3.5E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.050 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=1.100
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS BSIM4:
* low leakage
.MODEL P1 PMOS LEVEL=14 VTO=-0.45 U0=0.018 TOX= 3.5E-9 LINT=0.010U 
+K1 =0.450 K2=0.100 DVT0=2.300
+DVT1=0.540 LPE0=23.000e-9 ETA0=0.080
+NFACTOR=  1.6 U0=0.018 UA=3.000e-15
+WINT=0.020U LPE0=23.000e-9 
+KT1=-0.060 UTE=-1.800 VOFF=0.050
+XJ=0.150U NDEP=170.000e15 PCLM=0.700
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.30PS 50.00N
.PROBE
.END
